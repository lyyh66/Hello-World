module reg_test #
